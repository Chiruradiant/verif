module top;

initial 
$display("Hello World");

endmodule
