module top;

initial begin
$display("Hello World");
$display("Hi Eajaz");
end
endmodule
