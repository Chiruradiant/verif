module top;

initial begin
$display("Hello World");
$display("Hi Eajaz");
$display("Hi Gyani");
end
endmodule
